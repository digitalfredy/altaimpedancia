module Cero (/*AUTOARG*/
   // Outputs
   Salida
   ) ;
   output [15:0] Salida;

   assign Salida = 16'h0;
endmodule // Cero
